* STM32F103 Clock System Model - Super Simple Version
.SUBCKT STM32F103_CLOCK HSE VSS SYSCLK PLL_CLK HCLK PCLK1 PCLK2

* Simple RC buffers only - no flip-flops or complex logic
R1 HSE SYSCLK 10k
C1 SYSCLK VSS 100p

R2 SYSCLK PLL_CLK 10k
C2 PLL_CLK VSS 100p

R3 PLL_CLK HCLK 10k
C3 HCLK VSS 100p

R4 HCLK PCLK1 10k
C4 PCLK1 VSS 100p

R5 HCLK PCLK2 10k
C5 PCLK2 VSS 100p

.ENDS
